

module SAR_ADC_SVA /*#(
    parameter DATA_WIDTH = 32				 ,
    parameter ADDR_WIDTH = 32				 ,
    parameter NO_SLAVES  = 1					
) */(

input clk
);

endmodule : SAR_ADC_SVA